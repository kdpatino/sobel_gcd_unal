/home/dnmaldonador/Documents/sobel_gcd_unal/src/sobel_enhancement/src/verilog/sobel_core.sv