/home/dnmaldonador/Documents/sobel_gcd_unal/src/GCD/src/include/gcd.svh