/home/dnmaldonador/Documents/sobel_gcd_unal/src/spi_dep/verilog/spi_dep.sv