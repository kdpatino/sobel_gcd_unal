/home/dnmaldonador/Documents/sobel_gcd_unal/src/GCD/src/verilog/gcd_top.sv