/home/dnmaldonador/Documents/sobel_gcd_unal/src/spi_dep/verilog/adc_spi.sv